library ieee;
use ieee.std_logic_1164.all;

package globals is
    Constant N : integer := 32;
    constant M : integer := 2;
end;
